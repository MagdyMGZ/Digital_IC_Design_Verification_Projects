////////////////////////////////////////////////////////////////////////////////
// Author: Magdy Ahmed Abbas
// Company: Consultix 
// Description: Log2 Verilog Design
////////////////////////////////////////////////////////////////////////////////
module log2 #(
    parameter WIDTH = 32       // Q8.24 (8 bits for integer part + 24 bits for fraction part) to achieve error < 0.1 dB
) (
    input       wire        [WIDTH-1:0]      log2_in,       // 32 bit Integer Input
    input       wire                         clk,
    input       wire                         rstn,
    input       wire                         enable_in,
    output      reg                          valid_out,
    output      reg         [WIDTH-1:0]      log2_out       // log2_out[31:24] = Integer Part, log2_out[23:0] = Fraction Part
);

// log2(X) = N + log2(1 + F)
// N: integer part = position of MSB one in X
// F: fraction remainder after removing the MSB

reg [23:0] ROM [0:1023];

reg             enable_in_reg;
reg [WIDTH-1:0] log2_in_reg;
reg [WIDTH-1:0] log2_in_normalized;

reg [7:0]  int_part;
reg [23:0] frac_part;
reg [9:0]  frac_index;

// Register the Inputs
always @(posedge clk or negedge rstn) begin
    if (!rstn) begin
        enable_in_reg <= 0;
        log2_in_reg <= 0;
    end
    else if (enable_in) begin
        enable_in_reg <= enable_in;
        log2_in_reg <= log2_in;
    end
    else begin
        enable_in_reg <= 0;
        log2_in_reg <= 0;
    end
end

// Compute Integer and Fraction Parts
always @(*) begin
    if (enable_in_reg) begin
        int_part = log2_int(log2_in_reg);
        log2_in_normalized = log2_in_reg << (31 - int_part);
        frac_index = log2_in_normalized[30:21];        
        frac_part = ROM[frac_index];
    end
    else begin
        int_part = 0;
        frac_part = 0;
        frac_index = 0;
        log2_in_normalized = 0;
    end
end

// Output Block
always @(posedge clk or negedge rstn) begin
    if (!rstn) begin
        log2_out  <= 0;
        valid_out <= 0;
    end
    else if (enable_in_reg) begin
        log2_out <= {int_part,frac_part};
        valid_out <= 1;
    end
    else begin
        log2_out <= 0;
        valid_out <= 0;
    end
end

// LOD (Leading One Detector) Algorithm to get Most Significant One (Integer Part)
function reg [7:0] log2_int (input reg [31:0] value);
    integer i;
    reg flag;
    begin
        flag = 0;
        log2_int = 0;
        for (i = 31 ; i >= 0 ; i = i - 1) begin
            if (value[i] && !flag) begin
                log2_int = i;
                flag = 1;
            end
        end
    end
endfunction

// LUT (ROM) for log2(1 + k/1024) * 10000
always @(posedge clk or negedge rstn) begin
    if (!rstn) begin
        ROM[0] <= 0; ROM[1] <= 0; ROM[2] <= 0; ROM[3] <= 0; ROM[4] <= 0; ROM[5] <= 0; ROM[6] <= 0; ROM[7] <= 0; 
        ROM[8] <= 0; ROM[9] <= 0; ROM[10] <= 0; ROM[11] <= 0; ROM[12] <= 0; ROM[13] <= 0; ROM[14] <= 0; ROM[15] <= 0; 
        ROM[16] <= 0; ROM[17] <= 0; ROM[18] <= 0; ROM[19] <= 0; ROM[20] <= 0; ROM[21] <= 0; ROM[22] <= 0; ROM[23] <= 0; 
        ROM[24] <= 0; ROM[25] <= 0; ROM[26] <= 0; ROM[27] <= 0; ROM[28] <= 0; ROM[29] <= 0; ROM[30] <= 0; ROM[31] <= 0; 
        ROM[32] <= 0; ROM[33] <= 0; ROM[34] <= 0; ROM[35] <= 0; ROM[36] <= 0; ROM[37] <= 0; ROM[38] <= 0; ROM[39] <= 0; 
        ROM[40] <= 0; ROM[41] <= 0; ROM[42] <= 0; ROM[43] <= 0; ROM[44] <= 0; ROM[45] <= 0; ROM[46] <= 0; ROM[47] <= 0; 
        ROM[48] <= 0; ROM[49] <= 0; ROM[50] <= 0; ROM[51] <= 0; ROM[52] <= 0; ROM[53] <= 0; ROM[54] <= 0; ROM[55] <= 0; 
        ROM[56] <= 0; ROM[57] <= 0; ROM[58] <= 0; ROM[59] <= 0; ROM[60] <= 0; ROM[61] <= 0; ROM[62] <= 0; ROM[63] <= 0; 
        ROM[64] <= 0; ROM[65] <= 0; ROM[66] <= 0; ROM[67] <= 0; ROM[68] <= 0; ROM[69] <= 0; ROM[70] <= 0; ROM[71] <= 0; 
        ROM[72] <= 0; ROM[73] <= 0; ROM[74] <= 0; ROM[75] <= 0; ROM[76] <= 0; ROM[77] <= 0; ROM[78] <= 0; ROM[79] <= 0; 
        ROM[80] <= 0; ROM[81] <= 0; ROM[82] <= 0; ROM[83] <= 0; ROM[84] <= 0; ROM[85] <= 0; ROM[86] <= 0; ROM[87] <= 0; 
        ROM[88] <= 0; ROM[89] <= 0; ROM[90] <= 0; ROM[91] <= 0; ROM[92] <= 0; ROM[93] <= 0; ROM[94] <= 0; ROM[95] <= 0; 
        ROM[96] <= 0; ROM[97] <= 0; ROM[98] <= 0; ROM[99] <= 0; ROM[100] <= 0; ROM[101] <= 0; ROM[102] <= 0; ROM[103] <= 0; 
        ROM[104] <= 0; ROM[105] <= 0; ROM[106] <= 0; ROM[107] <= 0; ROM[108] <= 0; ROM[109] <= 0; ROM[110] <= 0; ROM[111] <= 0; 
        ROM[112] <= 0; ROM[113] <= 0; ROM[114] <= 0; ROM[115] <= 0; ROM[116] <= 0; ROM[117] <= 0; ROM[118] <= 0; ROM[119] <= 0; 
        ROM[120] <= 0; ROM[121] <= 0; ROM[122] <= 0; ROM[123] <= 0; ROM[124] <= 0; ROM[125] <= 0; ROM[126] <= 0; ROM[127] <= 0; 
        ROM[128] <= 0; ROM[129] <= 0; ROM[130] <= 0; ROM[131] <= 0; ROM[132] <= 0; ROM[133] <= 0; ROM[134] <= 0; ROM[135] <= 0; 
        ROM[136] <= 0; ROM[137] <= 0; ROM[138] <= 0; ROM[139] <= 0; ROM[140] <= 0; ROM[141] <= 0; ROM[142] <= 0; ROM[143] <= 0; 
        ROM[144] <= 0; ROM[145] <= 0; ROM[146] <= 0; ROM[147] <= 0; ROM[148] <= 0; ROM[149] <= 0; ROM[150] <= 0; ROM[151] <= 0; 
        ROM[152] <= 0; ROM[153] <= 0; ROM[154] <= 0; ROM[155] <= 0; ROM[156] <= 0; ROM[157] <= 0; ROM[158] <= 0; ROM[159] <= 0; 
        ROM[160] <= 0; ROM[161] <= 0; ROM[162] <= 0; ROM[163] <= 0; ROM[164] <= 0; ROM[165] <= 0; ROM[166] <= 0; ROM[167] <= 0; 
        ROM[168] <= 0; ROM[169] <= 0; ROM[170] <= 0; ROM[171] <= 0; ROM[172] <= 0; ROM[173] <= 0; ROM[174] <= 0; ROM[175] <= 0; 
        ROM[176] <= 0; ROM[177] <= 0; ROM[178] <= 0; ROM[179] <= 0; ROM[180] <= 0; ROM[181] <= 0; ROM[182] <= 0; ROM[183] <= 0; 
        ROM[184] <= 0; ROM[185] <= 0; ROM[186] <= 0; ROM[187] <= 0; ROM[188] <= 0; ROM[189] <= 0; ROM[190] <= 0; ROM[191] <= 0; 
        ROM[192] <= 0; ROM[193] <= 0; ROM[194] <= 0; ROM[195] <= 0; ROM[196] <= 0; ROM[197] <= 0; ROM[198] <= 0; ROM[199] <= 0; 
        ROM[200] <= 0; ROM[201] <= 0; ROM[202] <= 0; ROM[203] <= 0; ROM[204] <= 0; ROM[205] <= 0; ROM[206] <= 0; ROM[207] <= 0; 
        ROM[208] <= 0; ROM[209] <= 0; ROM[210] <= 0; ROM[211] <= 0; ROM[212] <= 0; ROM[213] <= 0; ROM[214] <= 0; ROM[215] <= 0; 
        ROM[216] <= 0; ROM[217] <= 0; ROM[218] <= 0; ROM[219] <= 0; ROM[220] <= 0; ROM[221] <= 0; ROM[222] <= 0; ROM[223] <= 0; 
        ROM[224] <= 0; ROM[225] <= 0; ROM[226] <= 0; ROM[227] <= 0; ROM[228] <= 0; ROM[229] <= 0; ROM[230] <= 0; ROM[231] <= 0; 
        ROM[232] <= 0; ROM[233] <= 0; ROM[234] <= 0; ROM[235] <= 0; ROM[236] <= 0; ROM[237] <= 0; ROM[238] <= 0; ROM[239] <= 0; 
        ROM[240] <= 0; ROM[241] <= 0; ROM[242] <= 0; ROM[243] <= 0; ROM[244] <= 0; ROM[245] <= 0; ROM[246] <= 0; ROM[247] <= 0; 
        ROM[248] <= 0; ROM[249] <= 0; ROM[250] <= 0; ROM[251] <= 0; ROM[252] <= 0; ROM[253] <= 0; ROM[254] <= 0; ROM[255] <= 0; 
        ROM[256] <= 0; ROM[257] <= 0; ROM[258] <= 0; ROM[259] <= 0; ROM[260] <= 0; ROM[261] <= 0; ROM[262] <= 0; ROM[263] <= 0; 
        ROM[264] <= 0; ROM[265] <= 0; ROM[266] <= 0; ROM[267] <= 0; ROM[268] <= 0; ROM[269] <= 0; ROM[270] <= 0; ROM[271] <= 0; 
        ROM[272] <= 0; ROM[273] <= 0; ROM[274] <= 0; ROM[275] <= 0; ROM[276] <= 0; ROM[277] <= 0; ROM[278] <= 0; ROM[279] <= 0; 
        ROM[280] <= 0; ROM[281] <= 0; ROM[282] <= 0; ROM[283] <= 0; ROM[284] <= 0; ROM[285] <= 0; ROM[286] <= 0; ROM[287] <= 0; 
        ROM[288] <= 0; ROM[289] <= 0; ROM[290] <= 0; ROM[291] <= 0; ROM[292] <= 0; ROM[293] <= 0; ROM[294] <= 0; ROM[295] <= 0; 
        ROM[296] <= 0; ROM[297] <= 0; ROM[298] <= 0; ROM[299] <= 0; ROM[300] <= 0; ROM[301] <= 0; ROM[302] <= 0; ROM[303] <= 0; 
        ROM[304] <= 0; ROM[305] <= 0; ROM[306] <= 0; ROM[307] <= 0; ROM[308] <= 0; ROM[309] <= 0; ROM[310] <= 0; ROM[311] <= 0; 
        ROM[312] <= 0; ROM[313] <= 0; ROM[314] <= 0; ROM[315] <= 0; ROM[316] <= 0; ROM[317] <= 0; ROM[318] <= 0; ROM[319] <= 0; 
        ROM[320] <= 0; ROM[321] <= 0; ROM[322] <= 0; ROM[323] <= 0; ROM[324] <= 0; ROM[325] <= 0; ROM[326] <= 0; ROM[327] <= 0; 
        ROM[328] <= 0; ROM[329] <= 0; ROM[330] <= 0; ROM[331] <= 0; ROM[332] <= 0; ROM[333] <= 0; ROM[334] <= 0; ROM[335] <= 0; 
        ROM[336] <= 0; ROM[337] <= 0; ROM[338] <= 0; ROM[339] <= 0; ROM[340] <= 0; ROM[341] <= 0; ROM[342] <= 0; ROM[343] <= 0; 
        ROM[344] <= 0; ROM[345] <= 0; ROM[346] <= 0; ROM[347] <= 0; ROM[348] <= 0; ROM[349] <= 0; ROM[350] <= 0; ROM[351] <= 0; 
        ROM[352] <= 0; ROM[353] <= 0; ROM[354] <= 0; ROM[355] <= 0; ROM[356] <= 0; ROM[357] <= 0; ROM[358] <= 0; ROM[359] <= 0; 
        ROM[360] <= 0; ROM[361] <= 0; ROM[362] <= 0; ROM[363] <= 0; ROM[364] <= 0; ROM[365] <= 0; ROM[366] <= 0; ROM[367] <= 0; 
        ROM[368] <= 0; ROM[369] <= 0; ROM[370] <= 0; ROM[371] <= 0; ROM[372] <= 0; ROM[373] <= 0; ROM[374] <= 0; ROM[375] <= 0; 
        ROM[376] <= 0; ROM[377] <= 0; ROM[378] <= 0; ROM[379] <= 0; ROM[380] <= 0; ROM[381] <= 0; ROM[382] <= 0; ROM[383] <= 0; 
        ROM[384] <= 0; ROM[385] <= 0; ROM[386] <= 0; ROM[387] <= 0; ROM[388] <= 0; ROM[389] <= 0; ROM[390] <= 0; ROM[391] <= 0; 
        ROM[392] <= 0; ROM[393] <= 0; ROM[394] <= 0; ROM[395] <= 0; ROM[396] <= 0; ROM[397] <= 0; ROM[398] <= 0; ROM[399] <= 0; 
        ROM[400] <= 0; ROM[401] <= 0; ROM[402] <= 0; ROM[403] <= 0; ROM[404] <= 0; ROM[405] <= 0; ROM[406] <= 0; ROM[407] <= 0; 
        ROM[408] <= 0; ROM[409] <= 0; ROM[410] <= 0; ROM[411] <= 0; ROM[412] <= 0; ROM[413] <= 0; ROM[414] <= 0; ROM[415] <= 0; 
        ROM[416] <= 0; ROM[417] <= 0; ROM[418] <= 0; ROM[419] <= 0; ROM[420] <= 0; ROM[421] <= 0; ROM[422] <= 0; ROM[423] <= 0; 
        ROM[424] <= 0; ROM[425] <= 0; ROM[426] <= 0; ROM[427] <= 0; ROM[428] <= 0; ROM[429] <= 0; ROM[430] <= 0; ROM[431] <= 0; 
        ROM[432] <= 0; ROM[433] <= 0; ROM[434] <= 0; ROM[435] <= 0; ROM[436] <= 0; ROM[437] <= 0; ROM[438] <= 0; ROM[439] <= 0; 
        ROM[440] <= 0; ROM[441] <= 0; ROM[442] <= 0; ROM[443] <= 0; ROM[444] <= 0; ROM[445] <= 0; ROM[446] <= 0; ROM[447] <= 0; 
        ROM[448] <= 0; ROM[449] <= 0; ROM[450] <= 0; ROM[451] <= 0; ROM[452] <= 0; ROM[453] <= 0; ROM[454] <= 0; ROM[455] <= 0; 
        ROM[456] <= 0; ROM[457] <= 0; ROM[458] <= 0; ROM[459] <= 0; ROM[460] <= 0; ROM[461] <= 0; ROM[462] <= 0; ROM[463] <= 0; 
        ROM[464] <= 0; ROM[465] <= 0; ROM[466] <= 0; ROM[467] <= 0; ROM[468] <= 0; ROM[469] <= 0; ROM[470] <= 0; ROM[471] <= 0; 
        ROM[472] <= 0; ROM[473] <= 0; ROM[474] <= 0; ROM[475] <= 0; ROM[476] <= 0; ROM[477] <= 0; ROM[478] <= 0; ROM[479] <= 0; 
        ROM[480] <= 0; ROM[481] <= 0; ROM[482] <= 0; ROM[483] <= 0; ROM[484] <= 0; ROM[485] <= 0; ROM[486] <= 0; ROM[487] <= 0; 
        ROM[488] <= 0; ROM[489] <= 0; ROM[490] <= 0; ROM[491] <= 0; ROM[492] <= 0; ROM[493] <= 0; ROM[494] <= 0; ROM[495] <= 0; 
        ROM[496] <= 0; ROM[497] <= 0; ROM[498] <= 0; ROM[499] <= 0; ROM[500] <= 0; ROM[501] <= 0; ROM[502] <= 0; ROM[503] <= 0; 
        ROM[504] <= 0; ROM[505] <= 0; ROM[506] <= 0; ROM[507] <= 0; ROM[508] <= 0; ROM[509] <= 0; ROM[510] <= 0; ROM[511] <= 0; 
        ROM[512] <= 0; ROM[513] <= 0; ROM[514] <= 0; ROM[515] <= 0; ROM[516] <= 0; ROM[517] <= 0; ROM[518] <= 0; ROM[519] <= 0; 
        ROM[520] <= 0; ROM[521] <= 0; ROM[522] <= 0; ROM[523] <= 0; ROM[524] <= 0; ROM[525] <= 0; ROM[526] <= 0; ROM[527] <= 0; 
        ROM[528] <= 0; ROM[529] <= 0; ROM[530] <= 0; ROM[531] <= 0; ROM[532] <= 0; ROM[533] <= 0; ROM[534] <= 0; ROM[535] <= 0; 
        ROM[536] <= 0; ROM[537] <= 0; ROM[538] <= 0; ROM[539] <= 0; ROM[540] <= 0; ROM[541] <= 0; ROM[542] <= 0; ROM[543] <= 0; 
        ROM[544] <= 0; ROM[545] <= 0; ROM[546] <= 0; ROM[547] <= 0; ROM[548] <= 0; ROM[549] <= 0; ROM[550] <= 0; ROM[551] <= 0; 
        ROM[552] <= 0; ROM[553] <= 0; ROM[554] <= 0; ROM[555] <= 0; ROM[556] <= 0; ROM[557] <= 0; ROM[558] <= 0; ROM[559] <= 0; 
        ROM[560] <= 0; ROM[561] <= 0; ROM[562] <= 0; ROM[563] <= 0; ROM[564] <= 0; ROM[565] <= 0; ROM[566] <= 0; ROM[567] <= 0; 
        ROM[568] <= 0; ROM[569] <= 0; ROM[570] <= 0; ROM[571] <= 0; ROM[572] <= 0; ROM[573] <= 0; ROM[574] <= 0; ROM[575] <= 0; 
        ROM[576] <= 0; ROM[577] <= 0; ROM[578] <= 0; ROM[579] <= 0; ROM[580] <= 0; ROM[581] <= 0; ROM[582] <= 0; ROM[583] <= 0; 
        ROM[584] <= 0; ROM[585] <= 0; ROM[586] <= 0; ROM[587] <= 0; ROM[588] <= 0; ROM[589] <= 0; ROM[590] <= 0; ROM[591] <= 0; 
        ROM[592] <= 0; ROM[593] <= 0; ROM[594] <= 0; ROM[595] <= 0; ROM[596] <= 0; ROM[597] <= 0; ROM[598] <= 0; ROM[599] <= 0; 
        ROM[600] <= 0; ROM[601] <= 0; ROM[602] <= 0; ROM[603] <= 0; ROM[604] <= 0; ROM[605] <= 0; ROM[606] <= 0; ROM[607] <= 0; 
        ROM[608] <= 0; ROM[609] <= 0; ROM[610] <= 0; ROM[611] <= 0; ROM[612] <= 0; ROM[613] <= 0; ROM[614] <= 0; ROM[615] <= 0; 
        ROM[616] <= 0; ROM[617] <= 0; ROM[618] <= 0; ROM[619] <= 0; ROM[620] <= 0; ROM[621] <= 0; ROM[622] <= 0; ROM[623] <= 0; 
        ROM[624] <= 0; ROM[625] <= 0; ROM[626] <= 0; ROM[627] <= 0; ROM[628] <= 0; ROM[629] <= 0; ROM[630] <= 0; ROM[631] <= 0; 
        ROM[632] <= 0; ROM[633] <= 0; ROM[634] <= 0; ROM[635] <= 0; ROM[636] <= 0; ROM[637] <= 0; ROM[638] <= 0; ROM[639] <= 0; 
        ROM[640] <= 0; ROM[641] <= 0; ROM[642] <= 0; ROM[643] <= 0; ROM[644] <= 0; ROM[645] <= 0; ROM[646] <= 0; ROM[647] <= 0; 
        ROM[648] <= 0; ROM[649] <= 0; ROM[650] <= 0; ROM[651] <= 0; ROM[652] <= 0; ROM[653] <= 0; ROM[654] <= 0; ROM[655] <= 0; 
        ROM[656] <= 0; ROM[657] <= 0; ROM[658] <= 0; ROM[659] <= 0; ROM[660] <= 0; ROM[661] <= 0; ROM[662] <= 0; ROM[663] <= 0; 
        ROM[664] <= 0; ROM[665] <= 0; ROM[666] <= 0; ROM[667] <= 0; ROM[668] <= 0; ROM[669] <= 0; ROM[670] <= 0; ROM[671] <= 0; 
        ROM[672] <= 0; ROM[673] <= 0; ROM[674] <= 0; ROM[675] <= 0; ROM[676] <= 0; ROM[677] <= 0; ROM[678] <= 0; ROM[679] <= 0; 
        ROM[680] <= 0; ROM[681] <= 0; ROM[682] <= 0; ROM[683] <= 0; ROM[684] <= 0; ROM[685] <= 0; ROM[686] <= 0; ROM[687] <= 0; 
        ROM[688] <= 0; ROM[689] <= 0; ROM[690] <= 0; ROM[691] <= 0; ROM[692] <= 0; ROM[693] <= 0; ROM[694] <= 0; ROM[695] <= 0; 
        ROM[696] <= 0; ROM[697] <= 0; ROM[698] <= 0; ROM[699] <= 0; ROM[700] <= 0; ROM[701] <= 0; ROM[702] <= 0; ROM[703] <= 0; 
        ROM[704] <= 0; ROM[705] <= 0; ROM[706] <= 0; ROM[707] <= 0; ROM[708] <= 0; ROM[709] <= 0; ROM[710] <= 0; ROM[711] <= 0; 
        ROM[712] <= 0; ROM[713] <= 0; ROM[714] <= 0; ROM[715] <= 0; ROM[716] <= 0; ROM[717] <= 0; ROM[718] <= 0; ROM[719] <= 0; 
        ROM[720] <= 0; ROM[721] <= 0; ROM[722] <= 0; ROM[723] <= 0; ROM[724] <= 0; ROM[725] <= 0; ROM[726] <= 0; ROM[727] <= 0; 
        ROM[728] <= 0; ROM[729] <= 0; ROM[730] <= 0; ROM[731] <= 0; ROM[732] <= 0; ROM[733] <= 0; ROM[734] <= 0; ROM[735] <= 0; 
        ROM[736] <= 0; ROM[737] <= 0; ROM[738] <= 0; ROM[739] <= 0; ROM[740] <= 0; ROM[741] <= 0; ROM[742] <= 0; ROM[743] <= 0; 
        ROM[744] <= 0; ROM[745] <= 0; ROM[746] <= 0; ROM[747] <= 0; ROM[748] <= 0; ROM[749] <= 0; ROM[750] <= 0; ROM[751] <= 0; 
        ROM[752] <= 0; ROM[753] <= 0; ROM[754] <= 0; ROM[755] <= 0; ROM[756] <= 0; ROM[757] <= 0; ROM[758] <= 0; ROM[759] <= 0; 
        ROM[760] <= 0; ROM[761] <= 0; ROM[762] <= 0; ROM[763] <= 0; ROM[764] <= 0; ROM[765] <= 0; ROM[766] <= 0; ROM[767] <= 0; 
        ROM[768] <= 0; ROM[769] <= 0; ROM[770] <= 0; ROM[771] <= 0; ROM[772] <= 0; ROM[773] <= 0; ROM[774] <= 0; ROM[775] <= 0; 
        ROM[776] <= 0; ROM[777] <= 0; ROM[778] <= 0; ROM[779] <= 0; ROM[780] <= 0; ROM[781] <= 0; ROM[782] <= 0; ROM[783] <= 0; 
        ROM[784] <= 0; ROM[785] <= 0; ROM[786] <= 0; ROM[787] <= 0; ROM[788] <= 0; ROM[789] <= 0; ROM[790] <= 0; ROM[791] <= 0; 
        ROM[792] <= 0; ROM[793] <= 0; ROM[794] <= 0; ROM[795] <= 0; ROM[796] <= 0; ROM[797] <= 0; ROM[798] <= 0; ROM[799] <= 0; 
        ROM[800] <= 0; ROM[801] <= 0; ROM[802] <= 0; ROM[803] <= 0; ROM[804] <= 0; ROM[805] <= 0; ROM[806] <= 0; ROM[807] <= 0; 
        ROM[808] <= 0; ROM[809] <= 0; ROM[810] <= 0; ROM[811] <= 0; ROM[812] <= 0; ROM[813] <= 0; ROM[814] <= 0; ROM[815] <= 0; 
        ROM[816] <= 0; ROM[817] <= 0; ROM[818] <= 0; ROM[819] <= 0; ROM[820] <= 0; ROM[821] <= 0; ROM[822] <= 0; ROM[823] <= 0; 
        ROM[824] <= 0; ROM[825] <= 0; ROM[826] <= 0; ROM[827] <= 0; ROM[828] <= 0; ROM[829] <= 0; ROM[830] <= 0; ROM[831] <= 0; 
        ROM[832] <= 0; ROM[833] <= 0; ROM[834] <= 0; ROM[835] <= 0; ROM[836] <= 0; ROM[837] <= 0; ROM[838] <= 0; ROM[839] <= 0; 
        ROM[840] <= 0; ROM[841] <= 0; ROM[842] <= 0; ROM[843] <= 0; ROM[844] <= 0; ROM[845] <= 0; ROM[846] <= 0; ROM[847] <= 0; 
        ROM[848] <= 0; ROM[849] <= 0; ROM[850] <= 0; ROM[851] <= 0; ROM[852] <= 0; ROM[853] <= 0; ROM[854] <= 0; ROM[855] <= 0; 
        ROM[856] <= 0; ROM[857] <= 0; ROM[858] <= 0; ROM[859] <= 0; ROM[860] <= 0; ROM[861] <= 0; ROM[862] <= 0; ROM[863] <= 0; 
        ROM[864] <= 0; ROM[865] <= 0; ROM[866] <= 0; ROM[867] <= 0; ROM[868] <= 0; ROM[869] <= 0; ROM[870] <= 0; ROM[871] <= 0; 
        ROM[872] <= 0; ROM[873] <= 0; ROM[874] <= 0; ROM[875] <= 0; ROM[876] <= 0; ROM[877] <= 0; ROM[878] <= 0; ROM[879] <= 0; 
        ROM[880] <= 0; ROM[881] <= 0; ROM[882] <= 0; ROM[883] <= 0; ROM[884] <= 0; ROM[885] <= 0; ROM[886] <= 0; ROM[887] <= 0; 
        ROM[888] <= 0; ROM[889] <= 0; ROM[890] <= 0; ROM[891] <= 0; ROM[892] <= 0; ROM[893] <= 0; ROM[894] <= 0; ROM[895] <= 0; 
        ROM[896] <= 0; ROM[897] <= 0; ROM[898] <= 0; ROM[899] <= 0; ROM[900] <= 0; ROM[901] <= 0; ROM[902] <= 0; ROM[903] <= 0; 
        ROM[904] <= 0; ROM[905] <= 0; ROM[906] <= 0; ROM[907] <= 0; ROM[908] <= 0; ROM[909] <= 0; ROM[910] <= 0; ROM[911] <= 0; 
        ROM[912] <= 0; ROM[913] <= 0; ROM[914] <= 0; ROM[915] <= 0; ROM[916] <= 0; ROM[917] <= 0; ROM[918] <= 0; ROM[919] <= 0; 
        ROM[920] <= 0; ROM[921] <= 0; ROM[922] <= 0; ROM[923] <= 0; ROM[924] <= 0; ROM[925] <= 0; ROM[926] <= 0; ROM[927] <= 0; 
        ROM[928] <= 0; ROM[929] <= 0; ROM[930] <= 0; ROM[931] <= 0; ROM[932] <= 0; ROM[933] <= 0; ROM[934] <= 0; ROM[935] <= 0; 
        ROM[936] <= 0; ROM[937] <= 0; ROM[938] <= 0; ROM[939] <= 0; ROM[940] <= 0; ROM[941] <= 0; ROM[942] <= 0; ROM[943] <= 0; 
        ROM[944] <= 0; ROM[945] <= 0; ROM[946] <= 0; ROM[947] <= 0; ROM[948] <= 0; ROM[949] <= 0; ROM[950] <= 0; ROM[951] <= 0; 
        ROM[952] <= 0; ROM[953] <= 0; ROM[954] <= 0; ROM[955] <= 0; ROM[956] <= 0; ROM[957] <= 0; ROM[958] <= 0; ROM[959] <= 0; 
        ROM[960] <= 0; ROM[961] <= 0; ROM[962] <= 0; ROM[963] <= 0; ROM[964] <= 0; ROM[965] <= 0; ROM[966] <= 0; ROM[967] <= 0; 
        ROM[968] <= 0; ROM[969] <= 0; ROM[970] <= 0; ROM[971] <= 0; ROM[972] <= 0; ROM[973] <= 0; ROM[974] <= 0; ROM[975] <= 0; 
        ROM[976] <= 0; ROM[977] <= 0; ROM[978] <= 0; ROM[979] <= 0; ROM[980] <= 0; ROM[981] <= 0; ROM[982] <= 0; ROM[983] <= 0; 
        ROM[984] <= 0; ROM[985] <= 0; ROM[986] <= 0; ROM[987] <= 0; ROM[988] <= 0; ROM[989] <= 0; ROM[990] <= 0; ROM[991] <= 0; 
        ROM[992] <= 0; ROM[993] <= 0; ROM[994] <= 0; ROM[995] <= 0; ROM[996] <= 0; ROM[997] <= 0; ROM[998] <= 0; ROM[999] <= 0; 
        ROM[1000] <= 0; ROM[1001] <= 0; ROM[1002] <= 0; ROM[1003] <= 0; ROM[1004] <= 0; ROM[1005] <= 0; ROM[1006] <= 0; ROM[1007] <= 0; 
        ROM[1008] <= 0; ROM[1009] <= 0; ROM[1010] <= 0; ROM[1011] <= 0; ROM[1012] <= 0; ROM[1013] <= 0; ROM[1014] <= 0; ROM[1015] <= 0; 
        ROM[1016] <= 0; ROM[1017] <= 0; ROM[1018] <= 0; ROM[1019] <= 0; ROM[1020] <= 0; ROM[1021] <= 0; ROM[1022] <= 0; ROM[1023] <= 0; 
    end
    else begin
        ROM[0] <= 24'd0; ROM[1] <= 24'd14; ROM[2] <= 24'd28; ROM[3] <= 24'd42; ROM[4] <= 24'd56; ROM[5] <= 24'd70; ROM[6] <= 24'd84; ROM[7] <= 24'd98; 
        ROM[8] <= 24'd112; ROM[9] <= 24'd126; ROM[10] <= 24'd140; ROM[11] <= 24'd154; ROM[12] <= 24'd168; ROM[13] <= 24'd182; ROM[14] <= 24'd196; ROM[15] <= 24'd210; 
        ROM[16] <= 24'd224; ROM[17] <= 24'd238; ROM[18] <= 24'd251; ROM[19] <= 24'd265; ROM[20] <= 24'd279; ROM[21] <= 24'd293; ROM[22] <= 24'd307; ROM[23] <= 24'd320; 
        ROM[24] <= 24'd334; ROM[25] <= 24'd348; ROM[26] <= 24'd362; ROM[27] <= 24'd375; ROM[28] <= 24'd389; ROM[29] <= 24'd403; ROM[30] <= 24'd417; ROM[31] <= 24'd430; 
        ROM[32] <= 24'd444; ROM[33] <= 24'd458; ROM[34] <= 24'd471; ROM[35] <= 24'd485; ROM[36] <= 24'd498; ROM[37] <= 24'd512; ROM[38] <= 24'd526; ROM[39] <= 24'd539; 
        ROM[40] <= 24'd553; ROM[41] <= 24'd566; ROM[42] <= 24'd580; ROM[43] <= 24'd593; ROM[44] <= 24'd607; ROM[45] <= 24'd620; ROM[46] <= 24'd634; ROM[47] <= 24'd647; 
        ROM[48] <= 24'd661; ROM[49] <= 24'd674; ROM[50] <= 24'd688; ROM[51] <= 24'd701; ROM[52] <= 24'd715; ROM[53] <= 24'd728; ROM[54] <= 24'd741; ROM[55] <= 24'd755; 
        ROM[56] <= 24'd768; ROM[57] <= 24'd782; ROM[58] <= 24'd795; ROM[59] <= 24'd808; ROM[60] <= 24'd821; ROM[61] <= 24'd835; ROM[62] <= 24'd848; ROM[63] <= 24'd861; 
        ROM[64] <= 24'd875; ROM[65] <= 24'd888; ROM[66] <= 24'd901; ROM[67] <= 24'd914; ROM[68] <= 24'd928; ROM[69] <= 24'd941; ROM[70] <= 24'd954; ROM[71] <= 24'd967; 
        ROM[72] <= 24'd980; ROM[73] <= 24'd993; ROM[74] <= 24'd1007; ROM[75] <= 24'd1020; ROM[76] <= 24'd1033; ROM[77] <= 24'd1046; ROM[78] <= 24'd1059; ROM[79] <= 24'd1072; 
        ROM[80] <= 24'd1085; ROM[81] <= 24'd1098; ROM[82] <= 24'd1111; ROM[83] <= 24'd1124; ROM[84] <= 24'd1137; ROM[85] <= 24'd1150; ROM[86] <= 24'd1163; ROM[87] <= 24'd1176; 
        ROM[88] <= 24'd1189; ROM[89] <= 24'd1202; ROM[90] <= 24'd1215; ROM[91] <= 24'd1228; ROM[92] <= 24'd1241; ROM[93] <= 24'd1254; ROM[94] <= 24'd1267; ROM[95] <= 24'd1280; 
        ROM[96] <= 24'd1293; ROM[97] <= 24'd1306; ROM[98] <= 24'd1319; ROM[99] <= 24'd1331; ROM[100] <= 24'd1344; ROM[101] <= 24'd1357; ROM[102] <= 24'd1370; ROM[103] <= 24'd1383; 
        ROM[104] <= 24'd1396; ROM[105] <= 24'd1408; ROM[106] <= 24'd1421; ROM[107] <= 24'd1434; ROM[108] <= 24'd1447; ROM[109] <= 24'd1459; ROM[110] <= 24'd1472; ROM[111] <= 24'd1485; 
        ROM[112] <= 24'd1497; ROM[113] <= 24'd1510; ROM[114] <= 24'd1523; ROM[115] <= 24'd1536; ROM[116] <= 24'd1548; ROM[117] <= 24'd1561; ROM[118] <= 24'd1573; ROM[119] <= 24'd1586; 
        ROM[120] <= 24'd1599; ROM[121] <= 24'd1611; ROM[122] <= 24'd1624; ROM[123] <= 24'd1636; ROM[124] <= 24'd1649; ROM[125] <= 24'd1662; ROM[126] <= 24'd1674; ROM[127] <= 24'd1687; 
        ROM[128] <= 24'd1699; ROM[129] <= 24'd1712; ROM[130] <= 24'd1724; ROM[131] <= 24'd1737; ROM[132] <= 24'd1749; ROM[133] <= 24'd1762; ROM[134] <= 24'd1774; ROM[135] <= 24'd1787; 
        ROM[136] <= 24'd1799; ROM[137] <= 24'd1812; ROM[138] <= 24'd1824; ROM[139] <= 24'd1836; ROM[140] <= 24'd1849; ROM[141] <= 24'd1861; ROM[142] <= 24'd1874; ROM[143] <= 24'd1886; 
        ROM[144] <= 24'd1898; ROM[145] <= 24'd1911; ROM[146] <= 24'd1923; ROM[147] <= 24'd1935; ROM[148] <= 24'd1948; ROM[149] <= 24'd1960; ROM[150] <= 24'd1972; ROM[151] <= 24'd1984; 
        ROM[152] <= 24'd1997; ROM[153] <= 24'd2009; ROM[154] <= 24'd2021; ROM[155] <= 24'd2033; ROM[156] <= 24'd2046; ROM[157] <= 24'd2058; ROM[158] <= 24'd2070; ROM[159] <= 24'd2082; 
        ROM[160] <= 24'd2095; ROM[161] <= 24'd2107; ROM[162] <= 24'd2119; ROM[163] <= 24'd2131; ROM[164] <= 24'd2143; ROM[165] <= 24'd2155; ROM[166] <= 24'd2167; ROM[167] <= 24'd2180; 
        ROM[168] <= 24'd2192; ROM[169] <= 24'd2204; ROM[170] <= 24'd2216; ROM[171] <= 24'd2228; ROM[172] <= 24'd2240; ROM[173] <= 24'd2252; ROM[174] <= 24'd2264; ROM[175] <= 24'd2276; 
        ROM[176] <= 24'd2288; ROM[177] <= 24'd2300; ROM[178] <= 24'd2312; ROM[179] <= 24'd2324; ROM[180] <= 24'd2336; ROM[181] <= 24'd2348; ROM[182] <= 24'd2360; ROM[183] <= 24'd2372; 
        ROM[184] <= 24'd2384; ROM[185] <= 24'd2396; ROM[186] <= 24'd2408; ROM[187] <= 24'd2420; ROM[188] <= 24'd2432; ROM[189] <= 24'd2444; ROM[190] <= 24'd2456; ROM[191] <= 24'd2467; 
        ROM[192] <= 24'd2479; ROM[193] <= 24'd2491; ROM[194] <= 24'd2503; ROM[195] <= 24'd2515; ROM[196] <= 24'd2527; ROM[197] <= 24'd2538; ROM[198] <= 24'd2550; ROM[199] <= 24'd2562; 
        ROM[200] <= 24'd2574; ROM[201] <= 24'd2586; ROM[202] <= 24'd2597; ROM[203] <= 24'd2609; ROM[204] <= 24'd2621; ROM[205] <= 24'd2633; ROM[206] <= 24'd2644; ROM[207] <= 24'd2656; 
        ROM[208] <= 24'd2668; ROM[209] <= 24'd2680; ROM[210] <= 24'd2691; ROM[211] <= 24'd2703; ROM[212] <= 24'd2715; ROM[213] <= 24'd2726; ROM[214] <= 24'd2738; ROM[215] <= 24'd2750; 
        ROM[216] <= 24'd2761; ROM[217] <= 24'd2773; ROM[218] <= 24'd2784; ROM[219] <= 24'd2796; ROM[220] <= 24'd2808; ROM[221] <= 24'd2819; ROM[222] <= 24'd2831; ROM[223] <= 24'd2842; 
        ROM[224] <= 24'd2854; ROM[225] <= 24'd2866; ROM[226] <= 24'd2877; ROM[227] <= 24'd2889; ROM[228] <= 24'd2900; ROM[229] <= 24'd2912; ROM[230] <= 24'd2923; ROM[231] <= 24'd2935; 
        ROM[232] <= 24'd2946; ROM[233] <= 24'd2958; ROM[234] <= 24'd2969; ROM[235] <= 24'd2981; ROM[236] <= 24'd2992; ROM[237] <= 24'd3004; ROM[238] <= 24'd3015; ROM[239] <= 24'd3026; 
        ROM[240] <= 24'd3038; ROM[241] <= 24'd3049; ROM[242] <= 24'd3061; ROM[243] <= 24'd3072; ROM[244] <= 24'd3083; ROM[245] <= 24'd3095; ROM[246] <= 24'd3106; ROM[247] <= 24'd3117; 
        ROM[248] <= 24'd3129; ROM[249] <= 24'd3140; ROM[250] <= 24'd3151; ROM[251] <= 24'd3163; ROM[252] <= 24'd3174; ROM[253] <= 24'd3185; ROM[254] <= 24'd3197; ROM[255] <= 24'd3208; 
        ROM[256] <= 24'd3219; ROM[257] <= 24'd3231; ROM[258] <= 24'd3242; ROM[259] <= 24'd3253; ROM[260] <= 24'd3264; ROM[261] <= 24'd3276; ROM[262] <= 24'd3287; ROM[263] <= 24'd3298; 
        ROM[264] <= 24'd3309; ROM[265] <= 24'd3320; ROM[266] <= 24'd3332; ROM[267] <= 24'd3343; ROM[268] <= 24'd3354; ROM[269] <= 24'd3365; ROM[270] <= 24'd3376; ROM[271] <= 24'd3387; 
        ROM[272] <= 24'd3399; ROM[273] <= 24'd3410; ROM[274] <= 24'd3421; ROM[275] <= 24'd3432; ROM[276] <= 24'd3443; ROM[277] <= 24'd3454; ROM[278] <= 24'd3465; ROM[279] <= 24'd3476; 
        ROM[280] <= 24'd3487; ROM[281] <= 24'd3498; ROM[282] <= 24'd3509; ROM[283] <= 24'd3520; ROM[284] <= 24'd3531; ROM[285] <= 24'd3542; ROM[286] <= 24'd3554; ROM[287] <= 24'd3565; 
        ROM[288] <= 24'd3576; ROM[289] <= 24'd3587; ROM[290] <= 24'd3597; ROM[291] <= 24'd3608; ROM[292] <= 24'd3619; ROM[293] <= 24'd3630; ROM[294] <= 24'd3641; ROM[295] <= 24'd3652; 
        ROM[296] <= 24'd3663; ROM[297] <= 24'd3674; ROM[298] <= 24'd3685; ROM[299] <= 24'd3696; ROM[300] <= 24'd3707; ROM[301] <= 24'd3718; ROM[302] <= 24'd3729; ROM[303] <= 24'd3740; 
        ROM[304] <= 24'd3750; ROM[305] <= 24'd3761; ROM[306] <= 24'd3772; ROM[307] <= 24'd3783; ROM[308] <= 24'd3794; ROM[309] <= 24'd3805; ROM[310] <= 24'd3815; ROM[311] <= 24'd3826; 
        ROM[312] <= 24'd3837; ROM[313] <= 24'd3848; ROM[314] <= 24'd3859; ROM[315] <= 24'd3869; ROM[316] <= 24'd3880; ROM[317] <= 24'd3891; ROM[318] <= 24'd3902; ROM[319] <= 24'd3912; 
        ROM[320] <= 24'd3923; ROM[321] <= 24'd3934; ROM[322] <= 24'd3945; ROM[323] <= 24'd3955; ROM[324] <= 24'd3966; ROM[325] <= 24'd3977; ROM[326] <= 24'd3987; ROM[327] <= 24'd3998; 
        ROM[328] <= 24'd4009; ROM[329] <= 24'd4019; ROM[330] <= 24'd4030; ROM[331] <= 24'd4041; ROM[332] <= 24'd4051; ROM[333] <= 24'd4062; ROM[334] <= 24'd4073; ROM[335] <= 24'd4083; 
        ROM[336] <= 24'd4094; ROM[337] <= 24'd4105; ROM[338] <= 24'd4115; ROM[339] <= 24'd4126; ROM[340] <= 24'd4136; ROM[341] <= 24'd4147; ROM[342] <= 24'd4157; ROM[343] <= 24'd4168; 
        ROM[344] <= 24'd4179; ROM[345] <= 24'd4189; ROM[346] <= 24'd4200; ROM[347] <= 24'd4210; ROM[348] <= 24'd4221; ROM[349] <= 24'd4231; ROM[350] <= 24'd4242; ROM[351] <= 24'd4252; 
        ROM[352] <= 24'd4263; ROM[353] <= 24'd4273; ROM[354] <= 24'd4284; ROM[355] <= 24'd4294; ROM[356] <= 24'd4305; ROM[357] <= 24'd4315; ROM[358] <= 24'd4325; ROM[359] <= 24'd4336; 
        ROM[360] <= 24'd4346; ROM[361] <= 24'd4357; ROM[362] <= 24'd4367; ROM[363] <= 24'd4378; ROM[364] <= 24'd4388; ROM[365] <= 24'd4398; ROM[366] <= 24'd4409; ROM[367] <= 24'd4419; 
        ROM[368] <= 24'd4429; ROM[369] <= 24'd4440; ROM[370] <= 24'd4450; ROM[371] <= 24'd4460; ROM[372] <= 24'd4471; ROM[373] <= 24'd4481; ROM[374] <= 24'd4491; ROM[375] <= 24'd4502; 
        ROM[376] <= 24'd4512; ROM[377] <= 24'd4522; ROM[378] <= 24'd4533; ROM[379] <= 24'd4543; ROM[380] <= 24'd4553; ROM[381] <= 24'd4564; ROM[382] <= 24'd4574; ROM[383] <= 24'd4584; 
        ROM[384] <= 24'd4594; ROM[385] <= 24'd4605; ROM[386] <= 24'd4615; ROM[387] <= 24'd4625; ROM[388] <= 24'd4635; ROM[389] <= 24'd4645; ROM[390] <= 24'd4656; ROM[391] <= 24'd4666; 
        ROM[392] <= 24'd4676; ROM[393] <= 24'd4686; ROM[394] <= 24'd4696; ROM[395] <= 24'd4707; ROM[396] <= 24'd4717; ROM[397] <= 24'd4727; ROM[398] <= 24'd4737; ROM[399] <= 24'd4747; 
        ROM[400] <= 24'd4757; ROM[401] <= 24'd4767; ROM[402] <= 24'd4778; ROM[403] <= 24'd4788; ROM[404] <= 24'd4798; ROM[405] <= 24'd4808; ROM[406] <= 24'd4818; ROM[407] <= 24'd4828; 
        ROM[408] <= 24'd4838; ROM[409] <= 24'd4848; ROM[410] <= 24'd4858; ROM[411] <= 24'd4868; ROM[412] <= 24'd4878; ROM[413] <= 24'd4888; ROM[414] <= 24'd4898; ROM[415] <= 24'd4909; 
        ROM[416] <= 24'd4919; ROM[417] <= 24'd4929; ROM[418] <= 24'd4939; ROM[419] <= 24'd4949; ROM[420] <= 24'd4959; ROM[421] <= 24'd4969; ROM[422] <= 24'd4979; ROM[423] <= 24'd4988; 
        ROM[424] <= 24'd4998; ROM[425] <= 24'd5008; ROM[426] <= 24'd5018; ROM[427] <= 24'd5028; ROM[428] <= 24'd5038; ROM[429] <= 24'd5048; ROM[430] <= 24'd5058; ROM[431] <= 24'd5068; 
        ROM[432] <= 24'd5078; ROM[433] <= 24'd5088; ROM[434] <= 24'd5098; ROM[435] <= 24'd5108; ROM[436] <= 24'd5118; ROM[437] <= 24'd5127; ROM[438] <= 24'd5137; ROM[439] <= 24'd5147; 
        ROM[440] <= 24'd5157; ROM[441] <= 24'd5167; ROM[442] <= 24'd5177; ROM[443] <= 24'd5187; ROM[444] <= 24'd5196; ROM[445] <= 24'd5206; ROM[446] <= 24'd5216; ROM[447] <= 24'd5226; 
        ROM[448] <= 24'd5236; ROM[449] <= 24'd5245; ROM[450] <= 24'd5255; ROM[451] <= 24'd5265; ROM[452] <= 24'd5275; ROM[453] <= 24'd5285; ROM[454] <= 24'd5294; ROM[455] <= 24'd5304; 
        ROM[456] <= 24'd5314; ROM[457] <= 24'd5324; ROM[458] <= 24'd5333; ROM[459] <= 24'd5343; ROM[460] <= 24'd5353; ROM[461] <= 24'd5362; ROM[462] <= 24'd5372; ROM[463] <= 24'd5382; 
        ROM[464] <= 24'd5392; ROM[465] <= 24'd5401; ROM[466] <= 24'd5411; ROM[467] <= 24'd5421; ROM[468] <= 24'd5430; ROM[469] <= 24'd5440; ROM[470] <= 24'd5450; ROM[471] <= 24'd5459; 
        ROM[472] <= 24'd5469; ROM[473] <= 24'd5479; ROM[474] <= 24'd5488; ROM[475] <= 24'd5498; ROM[476] <= 24'd5507; ROM[477] <= 24'd5517; ROM[478] <= 24'd5527; ROM[479] <= 24'd5536; 
        ROM[480] <= 24'd5546; ROM[481] <= 24'd5555; ROM[482] <= 24'd5565; ROM[483] <= 24'd5575; ROM[484] <= 24'd5584; ROM[485] <= 24'd5594; ROM[486] <= 24'd5603; ROM[487] <= 24'd5613; 
        ROM[488] <= 24'd5622; ROM[489] <= 24'd5632; ROM[490] <= 24'd5641; ROM[491] <= 24'd5651; ROM[492] <= 24'd5661; ROM[493] <= 24'd5670; ROM[494] <= 24'd5680; ROM[495] <= 24'd5689; 
        ROM[496] <= 24'd5699; ROM[497] <= 24'd5708; ROM[498] <= 24'd5718; ROM[499] <= 24'd5727; ROM[500] <= 24'd5736; ROM[501] <= 24'd5746; ROM[502] <= 24'd5755; ROM[503] <= 24'd5765; 
        ROM[504] <= 24'd5774; ROM[505] <= 24'd5784; ROM[506] <= 24'd5793; ROM[507] <= 24'd5803; ROM[508] <= 24'd5812; ROM[509] <= 24'd5821; ROM[510] <= 24'd5831; ROM[511] <= 24'd5840; 
        ROM[512] <= 24'd5850; ROM[513] <= 24'd5859; ROM[514] <= 24'd5868; ROM[515] <= 24'd5878; ROM[516] <= 24'd5887; ROM[517] <= 24'd5897; ROM[518] <= 24'd5906; ROM[519] <= 24'd5915; 
        ROM[520] <= 24'd5925; ROM[521] <= 24'd5934; ROM[522] <= 24'd5943; ROM[523] <= 24'd5953; ROM[524] <= 24'd5962; ROM[525] <= 24'd5971; ROM[526] <= 24'd5981; ROM[527] <= 24'd5990; 
        ROM[528] <= 24'd5999; ROM[529] <= 24'd6008; ROM[530] <= 24'd6018; ROM[531] <= 24'd6027; ROM[532] <= 24'd6036; ROM[533] <= 24'd6046; ROM[534] <= 24'd6055; ROM[535] <= 24'd6064; 
        ROM[536] <= 24'd6073; ROM[537] <= 24'd6083; ROM[538] <= 24'd6092; ROM[539] <= 24'd6101; ROM[540] <= 24'd6110; ROM[541] <= 24'd6119; ROM[542] <= 24'd6129; ROM[543] <= 24'd6138; 
        ROM[544] <= 24'd6147; ROM[545] <= 24'd6156; ROM[546] <= 24'd6165; ROM[547] <= 24'd6175; ROM[548] <= 24'd6184; ROM[549] <= 24'd6193; ROM[550] <= 24'd6202; ROM[551] <= 24'd6211; 
        ROM[552] <= 24'd6221; ROM[553] <= 24'd6230; ROM[554] <= 24'd6239; ROM[555] <= 24'd6248; ROM[556] <= 24'd6257; ROM[557] <= 24'd6266; ROM[558] <= 24'd6275; ROM[559] <= 24'd6284; 
        ROM[560] <= 24'd6294; ROM[561] <= 24'd6303; ROM[562] <= 24'd6312; ROM[563] <= 24'd6321; ROM[564] <= 24'd6330; ROM[565] <= 24'd6339; ROM[566] <= 24'd6348; ROM[567] <= 24'd6357; 
        ROM[568] <= 24'd6366; ROM[569] <= 24'd6375; ROM[570] <= 24'd6384; ROM[571] <= 24'd6393; ROM[572] <= 24'd6402; ROM[573] <= 24'd6411; ROM[574] <= 24'd6421; ROM[575] <= 24'd6430; 
        ROM[576] <= 24'd6439; ROM[577] <= 24'd6448; ROM[578] <= 24'd6457; ROM[579] <= 24'd6466; ROM[580] <= 24'd6475; ROM[581] <= 24'd6484; ROM[582] <= 24'd6493; ROM[583] <= 24'd6502; 
        ROM[584] <= 24'd6511; ROM[585] <= 24'd6519; ROM[586] <= 24'd6528; ROM[587] <= 24'd6537; ROM[588] <= 24'd6546; ROM[589] <= 24'd6555; ROM[590] <= 24'd6564; ROM[591] <= 24'd6573; 
        ROM[592] <= 24'd6582; ROM[593] <= 24'd6591; ROM[594] <= 24'd6600; ROM[595] <= 24'd6609; ROM[596] <= 24'd6618; ROM[597] <= 24'd6627; ROM[598] <= 24'd6636; ROM[599] <= 24'd6644; 
        ROM[600] <= 24'd6653; ROM[601] <= 24'd6662; ROM[602] <= 24'd6671; ROM[603] <= 24'd6680; ROM[604] <= 24'd6689; ROM[605] <= 24'd6698; ROM[606] <= 24'd6707; ROM[607] <= 24'd6715; 
        ROM[608] <= 24'd6724; ROM[609] <= 24'd6733; ROM[610] <= 24'd6742; ROM[611] <= 24'd6751; ROM[612] <= 24'd6760; ROM[613] <= 24'd6768; ROM[614] <= 24'd6777; ROM[615] <= 24'd6786; 
        ROM[616] <= 24'd6795; ROM[617] <= 24'd6804; ROM[618] <= 24'd6812; ROM[619] <= 24'd6821; ROM[620] <= 24'd6830; ROM[621] <= 24'd6839; ROM[622] <= 24'd6847; ROM[623] <= 24'd6856; 
        ROM[624] <= 24'd6865; ROM[625] <= 24'd6874; ROM[626] <= 24'd6883; ROM[627] <= 24'd6891; ROM[628] <= 24'd6900; ROM[629] <= 24'd6909; ROM[630] <= 24'd6917; ROM[631] <= 24'd6926; 
        ROM[632] <= 24'd6935; ROM[633] <= 24'd6944; ROM[634] <= 24'd6952; ROM[635] <= 24'd6961; ROM[636] <= 24'd6970; ROM[637] <= 24'd6978; ROM[638] <= 24'd6987; ROM[639] <= 24'd6996; 
        ROM[640] <= 24'd7004; ROM[641] <= 24'd7013; ROM[642] <= 24'd7022; ROM[643] <= 24'd7030; ROM[644] <= 24'd7039; ROM[645] <= 24'd7048; ROM[646] <= 24'd7056; ROM[647] <= 24'd7065; 
        ROM[648] <= 24'd7074; ROM[649] <= 24'd7082; ROM[650] <= 24'd7091; ROM[651] <= 24'd7099; ROM[652] <= 24'd7108; ROM[653] <= 24'd7117; ROM[654] <= 24'd7125; ROM[655] <= 24'd7134; 
        ROM[656] <= 24'd7142; ROM[657] <= 24'd7151; ROM[658] <= 24'd7160; ROM[659] <= 24'd7168; ROM[660] <= 24'd7177; ROM[661] <= 24'd7185; ROM[662] <= 24'd7194; ROM[663] <= 24'd7202; 
        ROM[664] <= 24'd7211; ROM[665] <= 24'd7220; ROM[666] <= 24'd7228; ROM[667] <= 24'd7237; ROM[668] <= 24'd7245; ROM[669] <= 24'd7254; ROM[670] <= 24'd7262; ROM[671] <= 24'd7271; 
        ROM[672] <= 24'd7279; ROM[673] <= 24'd7288; ROM[674] <= 24'd7296; ROM[675] <= 24'd7305; ROM[676] <= 24'd7313; ROM[677] <= 24'd7322; ROM[678] <= 24'd7330; ROM[679] <= 24'd7339; 
        ROM[680] <= 24'd7347; ROM[681] <= 24'd7356; ROM[682] <= 24'd7364; ROM[683] <= 24'd7372; ROM[684] <= 24'd7381; ROM[685] <= 24'd7389; ROM[686] <= 24'd7398; ROM[687] <= 24'd7406; 
        ROM[688] <= 24'd7415; ROM[689] <= 24'd7423; ROM[690] <= 24'd7432; ROM[691] <= 24'd7440; ROM[692] <= 24'd7448; ROM[693] <= 24'd7457; ROM[694] <= 24'd7465; ROM[695] <= 24'd7474; 
        ROM[696] <= 24'd7482; ROM[697] <= 24'd7490; ROM[698] <= 24'd7499; ROM[699] <= 24'd7507; ROM[700] <= 24'd7515; ROM[701] <= 24'd7524; ROM[702] <= 24'd7532; ROM[703] <= 24'd7541; 
        ROM[704] <= 24'd7549; ROM[705] <= 24'd7557; ROM[706] <= 24'd7566; ROM[707] <= 24'd7574; ROM[708] <= 24'd7582; ROM[709] <= 24'd7591; ROM[710] <= 24'd7599; ROM[711] <= 24'd7607; 
        ROM[712] <= 24'd7616; ROM[713] <= 24'd7624; ROM[714] <= 24'd7632; ROM[715] <= 24'd7640; ROM[716] <= 24'd7649; ROM[717] <= 24'd7657; ROM[718] <= 24'd7665; ROM[719] <= 24'd7674; 
        ROM[720] <= 24'd7682; ROM[721] <= 24'd7690; ROM[722] <= 24'd7698; ROM[723] <= 24'd7707; ROM[724] <= 24'd7715; ROM[725] <= 24'd7723; ROM[726] <= 24'd7731; ROM[727] <= 24'd7740; 
        ROM[728] <= 24'd7748; ROM[729] <= 24'd7756; ROM[730] <= 24'd7764; ROM[731] <= 24'd7773; ROM[732] <= 24'd7781; ROM[733] <= 24'd7789; ROM[734] <= 24'd7797; ROM[735] <= 24'd7805; 
        ROM[736] <= 24'd7814; ROM[737] <= 24'd7822; ROM[738] <= 24'd7830; ROM[739] <= 24'd7838; ROM[740] <= 24'd7846; ROM[741] <= 24'd7855; ROM[742] <= 24'd7863; ROM[743] <= 24'd7871; 
        ROM[744] <= 24'd7879; ROM[745] <= 24'd7887; ROM[746] <= 24'd7895; ROM[747] <= 24'd7903; ROM[748] <= 24'd7912; ROM[749] <= 24'd7920; ROM[750] <= 24'd7928; ROM[751] <= 24'd7936; 
        ROM[752] <= 24'd7944; ROM[753] <= 24'd7952; ROM[754] <= 24'd7960; ROM[755] <= 24'd7969; ROM[756] <= 24'd7977; ROM[757] <= 24'd7985; ROM[758] <= 24'd7993; ROM[759] <= 24'd8001; 
        ROM[760] <= 24'd8009; ROM[761] <= 24'd8017; ROM[762] <= 24'd8025; ROM[763] <= 24'd8033; ROM[764] <= 24'd8041; ROM[765] <= 24'd8049; ROM[766] <= 24'd8057; ROM[767] <= 24'd8065; 
        ROM[768] <= 24'd8074; ROM[769] <= 24'd8082; ROM[770] <= 24'd8090; ROM[771] <= 24'd8098; ROM[772] <= 24'd8106; ROM[773] <= 24'd8114; ROM[774] <= 24'd8122; ROM[775] <= 24'd8130; 
        ROM[776] <= 24'd8138; ROM[777] <= 24'd8146; ROM[778] <= 24'd8154; ROM[779] <= 24'd8162; ROM[780] <= 24'd8170; ROM[781] <= 24'd8178; ROM[782] <= 24'd8186; ROM[783] <= 24'd8194; 
        ROM[784] <= 24'd8202; ROM[785] <= 24'd8210; ROM[786] <= 24'd8218; ROM[787] <= 24'd8226; ROM[788] <= 24'd8234; ROM[789] <= 24'd8242; ROM[790] <= 24'd8250; ROM[791] <= 24'd8258; 
        ROM[792] <= 24'd8265; ROM[793] <= 24'd8273; ROM[794] <= 24'd8281; ROM[795] <= 24'd8289; ROM[796] <= 24'd8297; ROM[797] <= 24'd8305; ROM[798] <= 24'd8313; ROM[799] <= 24'd8321; 
        ROM[800] <= 24'd8329; ROM[801] <= 24'd8337; ROM[802] <= 24'd8345; ROM[803] <= 24'd8353; ROM[804] <= 24'd8361; ROM[805] <= 24'd8368; ROM[806] <= 24'd8376; ROM[807] <= 24'd8384; 
        ROM[808] <= 24'd8392; ROM[809] <= 24'd8400; ROM[810] <= 24'd8408; ROM[811] <= 24'd8416; ROM[812] <= 24'd8424; ROM[813] <= 24'd8431; ROM[814] <= 24'd8439; ROM[815] <= 24'd8447; 
        ROM[816] <= 24'd8455; ROM[817] <= 24'd8463; ROM[818] <= 24'd8471; ROM[819] <= 24'd8478; ROM[820] <= 24'd8486; ROM[821] <= 24'd8494; ROM[822] <= 24'd8502; ROM[823] <= 24'd8510; 
        ROM[824] <= 24'd8517; ROM[825] <= 24'd8525; ROM[826] <= 24'd8533; ROM[827] <= 24'd8541; ROM[828] <= 24'd8549; ROM[829] <= 24'd8556; ROM[830] <= 24'd8564; ROM[831] <= 24'd8572; 
        ROM[832] <= 24'd8580; ROM[833] <= 24'd8588; ROM[834] <= 24'd8595; ROM[835] <= 24'd8603; ROM[836] <= 24'd8611; ROM[837] <= 24'd8619; ROM[838] <= 24'd8626; ROM[839] <= 24'd8634; 
        ROM[840] <= 24'd8642; ROM[841] <= 24'd8650; ROM[842] <= 24'd8657; ROM[843] <= 24'd8665; ROM[844] <= 24'd8673; ROM[845] <= 24'd8681; ROM[846] <= 24'd8688; ROM[847] <= 24'd8696; 
        ROM[848] <= 24'd8704; ROM[849] <= 24'd8711; ROM[850] <= 24'd8719; ROM[851] <= 24'd8727; ROM[852] <= 24'd8734; ROM[853] <= 24'd8742; ROM[854] <= 24'd8750; ROM[855] <= 24'd8757; 
        ROM[856] <= 24'd8765; ROM[857] <= 24'd8773; ROM[858] <= 24'd8781; ROM[859] <= 24'd8788; ROM[860] <= 24'd8796; ROM[861] <= 24'd8803; ROM[862] <= 24'd8811; ROM[863] <= 24'd8819; 
        ROM[864] <= 24'd8826; ROM[865] <= 24'd8834; ROM[866] <= 24'd8842; ROM[867] <= 24'd8849; ROM[868] <= 24'd8857; ROM[869] <= 24'd8865; ROM[870] <= 24'd8872; ROM[871] <= 24'd8880; 
        ROM[872] <= 24'd8887; ROM[873] <= 24'd8895; ROM[874] <= 24'd8903; ROM[875] <= 24'd8910; ROM[876] <= 24'd8918; ROM[877] <= 24'd8925; ROM[878] <= 24'd8933; ROM[879] <= 24'd8941; 
        ROM[880] <= 24'd8948; ROM[881] <= 24'd8956; ROM[882] <= 24'd8963; ROM[883] <= 24'd8971; ROM[884] <= 24'd8978; ROM[885] <= 24'd8986; ROM[886] <= 24'd8994; ROM[887] <= 24'd9001; 
        ROM[888] <= 24'd9009; ROM[889] <= 24'd9016; ROM[890] <= 24'd9024; ROM[891] <= 24'd9031; ROM[892] <= 24'd9039; ROM[893] <= 24'd9046; ROM[894] <= 24'd9054; ROM[895] <= 24'd9061; 
        ROM[896] <= 24'd9069; ROM[897] <= 24'd9076; ROM[898] <= 24'd9084; ROM[899] <= 24'd9091; ROM[900] <= 24'd9099; ROM[901] <= 24'd9106; ROM[902] <= 24'd9114; ROM[903] <= 24'd9121; 
        ROM[904] <= 24'd9129; ROM[905] <= 24'd9136; ROM[906] <= 24'd9144; ROM[907] <= 24'd9151; ROM[908] <= 24'd9159; ROM[909] <= 24'd9166; ROM[910] <= 24'd9174; ROM[911] <= 24'd9181; 
        ROM[912] <= 24'd9189; ROM[913] <= 24'd9196; ROM[914] <= 24'd9204; ROM[915] <= 24'd9211; ROM[916] <= 24'd9218; ROM[917] <= 24'd9226; ROM[918] <= 24'd9233; ROM[919] <= 24'd9241; 
        ROM[920] <= 24'd9248; ROM[921] <= 24'd9256; ROM[922] <= 24'd9263; ROM[923] <= 24'd9270; ROM[924] <= 24'd9278; ROM[925] <= 24'd9285; ROM[926] <= 24'd9293; ROM[927] <= 24'd9300; 
        ROM[928] <= 24'd9307; ROM[929] <= 24'd9315; ROM[930] <= 24'd9322; ROM[931] <= 24'd9330; ROM[932] <= 24'd9337; ROM[933] <= 24'd9344; ROM[934] <= 24'd9352; ROM[935] <= 24'd9359; 
        ROM[936] <= 24'd9366; ROM[937] <= 24'd9374; ROM[938] <= 24'd9381; ROM[939] <= 24'd9388; ROM[940] <= 24'd9396; ROM[941] <= 24'd9403; ROM[942] <= 24'd9410; ROM[943] <= 24'd9418; 
        ROM[944] <= 24'd9425; ROM[945] <= 24'd9432; ROM[946] <= 24'd9440; ROM[947] <= 24'd9447; ROM[948] <= 24'd9454; ROM[949] <= 24'd9462; ROM[950] <= 24'd9469; ROM[951] <= 24'd9476; 
        ROM[952] <= 24'd9484; ROM[953] <= 24'd9491; ROM[954] <= 24'd9498; ROM[955] <= 24'd9506; ROM[956] <= 24'd9513; ROM[957] <= 24'd9520; ROM[958] <= 24'd9527; ROM[959] <= 24'd9535; 
        ROM[960] <= 24'd9542; ROM[961] <= 24'd9549; ROM[962] <= 24'd9556; ROM[963] <= 24'd9564; ROM[964] <= 24'd9571; ROM[965] <= 24'd9578; ROM[966] <= 24'd9586; ROM[967] <= 24'd9593; 
        ROM[968] <= 24'd9600; ROM[969] <= 24'd9607; ROM[970] <= 24'd9614; ROM[971] <= 24'd9622; ROM[972] <= 24'd9629; ROM[973] <= 24'd9636; ROM[974] <= 24'd9643; ROM[975] <= 24'd9651; 
        ROM[976] <= 24'd9658; ROM[977] <= 24'd9665; ROM[978] <= 24'd9672; ROM[979] <= 24'd9679; ROM[980] <= 24'd9687; ROM[981] <= 24'd9694; ROM[982] <= 24'd9701; ROM[983] <= 24'd9708; 
        ROM[984] <= 24'd9715; ROM[985] <= 24'd9723; ROM[986] <= 24'd9730; ROM[987] <= 24'd9737; ROM[988] <= 24'd9744; ROM[989] <= 24'd9751; ROM[990] <= 24'd9758; ROM[991] <= 24'd9766; 
        ROM[992] <= 24'd9773; ROM[993] <= 24'd9780; ROM[994] <= 24'd9787; ROM[995] <= 24'd9794; ROM[996] <= 24'd9801; ROM[997] <= 24'd9809; ROM[998] <= 24'd9816; ROM[999] <= 24'd9823; 
        ROM[1000] <= 24'd9830; ROM[1001] <= 24'd9837; ROM[1002] <= 24'd9844; ROM[1003] <= 24'd9851; ROM[1004] <= 24'd9858; ROM[1005] <= 24'd9866; ROM[1006] <= 24'd9873; ROM[1007] <= 24'd9880; 
        ROM[1008] <= 24'd9887; ROM[1009] <= 24'd9894; ROM[1010] <= 24'd9901; ROM[1011] <= 24'd9908; ROM[1012] <= 24'd9915; ROM[1013] <= 24'd9922; ROM[1014] <= 24'd9929; ROM[1015] <= 24'd9936; 
        ROM[1016] <= 24'd9944; ROM[1017] <= 24'd9951; ROM[1018] <= 24'd9958; ROM[1019] <= 24'd9965; ROM[1020] <= 24'd9972; ROM[1021] <= 24'd9979; ROM[1022] <= 24'd9986; ROM[1023] <= 24'd9993; 
    end
end

endmodule

// localparam reg [23:0] ROM [0:1023] = '{
//     24'd0       , 24'd14      , 24'd28      , 24'd42      , 24'd56      , 24'd70      , 24'd84      , 24'd98      , 
//     24'd112     , 24'd126     , 24'd140     , 24'd154     , 24'd168     , 24'd182     , 24'd196     , 24'd210     , 
//     24'd224     , 24'd238     , 24'd251     , 24'd265     , 24'd279     , 24'd293     , 24'd307     , 24'd320     , 
//     24'd334     , 24'd348     , 24'd362     , 24'd375     , 24'd389     , 24'd403     , 24'd417     , 24'd430     , 
//     24'd444     , 24'd458     , 24'd471     , 24'd485     , 24'd498     , 24'd512     , 24'd526     , 24'd539     , 
//     24'd553     , 24'd566     , 24'd580     , 24'd593     , 24'd607     , 24'd620     , 24'd634     , 24'd647     , 
//     24'd661     , 24'd674     , 24'd688     , 24'd701     , 24'd715     , 24'd728     , 24'd741     , 24'd755     , 
//     24'd768     , 24'd782     , 24'd795     , 24'd808     , 24'd821     , 24'd835     , 24'd848     , 24'd861     , 
//     24'd875     , 24'd888     , 24'd901     , 24'd914     , 24'd928     , 24'd941     , 24'd954     , 24'd967     , 
//     24'd980     , 24'd993     , 24'd1007    , 24'd1020    , 24'd1033    , 24'd1046    , 24'd1059    , 24'd1072    , 
//     24'd1085    , 24'd1098    , 24'd1111    , 24'd1124    , 24'd1137    , 24'd1150    , 24'd1163    , 24'd1176    , 
//     24'd1189    , 24'd1202    , 24'd1215    , 24'd1228    , 24'd1241    , 24'd1254    , 24'd1267    , 24'd1280    , 
//     24'd1293    , 24'd1306    , 24'd1319    , 24'd1331    , 24'd1344    , 24'd1357    , 24'd1370    , 24'd1383    , 
//     24'd1396    , 24'd1408    , 24'd1421    , 24'd1434    , 24'd1447    , 24'd1459    , 24'd1472    , 24'd1485    , 
//     24'd1497    , 24'd1510    , 24'd1523    , 24'd1536    , 24'd1548    , 24'd1561    , 24'd1573    , 24'd1586    , 
//     24'd1599    , 24'd1611    , 24'd1624    , 24'd1636    , 24'd1649    , 24'd1662    , 24'd1674    , 24'd1687    , 
//     24'd1699    , 24'd1712    , 24'd1724    , 24'd1737    , 24'd1749    , 24'd1762    , 24'd1774    , 24'd1787    , 
//     24'd1799    , 24'd1812    , 24'd1824    , 24'd1836    , 24'd1849    , 24'd1861    , 24'd1874    , 24'd1886    , 
//     24'd1898    , 24'd1911    , 24'd1923    , 24'd1935    , 24'd1948    , 24'd1960    , 24'd1972    , 24'd1984    , 
//     24'd1997    , 24'd2009    , 24'd2021    , 24'd2033    , 24'd2046    , 24'd2058    , 24'd2070    , 24'd2082    , 
//     24'd2095    , 24'd2107    , 24'd2119    , 24'd2131    , 24'd2143    , 24'd2155    , 24'd2167    , 24'd2180    , 
//     24'd2192    , 24'd2204    , 24'd2216    , 24'd2228    , 24'd2240    , 24'd2252    , 24'd2264    , 24'd2276    , 
//     24'd2288    , 24'd2300    , 24'd2312    , 24'd2324    , 24'd2336    , 24'd2348    , 24'd2360    , 24'd2372    , 
//     24'd2384    , 24'd2396    , 24'd2408    , 24'd2420    , 24'd2432    , 24'd2444    , 24'd2456    , 24'd2467    , 
//     24'd2479    , 24'd2491    , 24'd2503    , 24'd2515    , 24'd2527    , 24'd2538    , 24'd2550    , 24'd2562    , 
//     24'd2574    , 24'd2586    , 24'd2597    , 24'd2609    , 24'd2621    , 24'd2633    , 24'd2644    , 24'd2656    , 
//     24'd2668    , 24'd2680    , 24'd2691    , 24'd2703    , 24'd2715    , 24'd2726    , 24'd2738    , 24'd2750    , 
//     24'd2761    , 24'd2773    , 24'd2784    , 24'd2796    , 24'd2808    , 24'd2819    , 24'd2831    , 24'd2842    , 
//     24'd2854    , 24'd2866    , 24'd2877    , 24'd2889    , 24'd2900    , 24'd2912    , 24'd2923    , 24'd2935    , 
//     24'd2946    , 24'd2958    , 24'd2969    , 24'd2981    , 24'd2992    , 24'd3004    , 24'd3015    , 24'd3026    , 
//     24'd3038    , 24'd3049    , 24'd3061    , 24'd3072    , 24'd3083    , 24'd3095    , 24'd3106    , 24'd3117    , 
//     24'd3129    , 24'd3140    , 24'd3151    , 24'd3163    , 24'd3174    , 24'd3185    , 24'd3197    , 24'd3208    , 
//     24'd3219    , 24'd3231    , 24'd3242    , 24'd3253    , 24'd3264    , 24'd3276    , 24'd3287    , 24'd3298    , 
//     24'd3309    , 24'd3320    , 24'd3332    , 24'd3343    , 24'd3354    , 24'd3365    , 24'd3376    , 24'd3387    , 
//     24'd3399    , 24'd3410    , 24'd3421    , 24'd3432    , 24'd3443    , 24'd3454    , 24'd3465    , 24'd3476    , 
//     24'd3487    , 24'd3498    , 24'd3509    , 24'd3520    , 24'd3531    , 24'd3542    , 24'd3554    , 24'd3565    , 
//     24'd3576    , 24'd3587    , 24'd3597    , 24'd3608    , 24'd3619    , 24'd3630    , 24'd3641    , 24'd3652    , 
//     24'd3663    , 24'd3674    , 24'd3685    , 24'd3696    , 24'd3707    , 24'd3718    , 24'd3729    , 24'd3740    , 
//     24'd3750    , 24'd3761    , 24'd3772    , 24'd3783    , 24'd3794    , 24'd3805    , 24'd3815    , 24'd3826    , 
//     24'd3837    , 24'd3848    , 24'd3859    , 24'd3869    , 24'd3880    , 24'd3891    , 24'd3902    , 24'd3912    , 
//     24'd3923    , 24'd3934    , 24'd3945    , 24'd3955    , 24'd3966    , 24'd3977    , 24'd3987    , 24'd3998    , 
//     24'd4009    , 24'd4019    , 24'd4030    , 24'd4041    , 24'd4051    , 24'd4062    , 24'd4073    , 24'd4083    , 
//     24'd4094    , 24'd4105    , 24'd4115    , 24'd4126    , 24'd4136    , 24'd4147    , 24'd4157    , 24'd4168    , 
//     24'd4179    , 24'd4189    , 24'd4200    , 24'd4210    , 24'd4221    , 24'd4231    , 24'd4242    , 24'd4252    , 
//     24'd4263    , 24'd4273    , 24'd4284    , 24'd4294    , 24'd4305    , 24'd4315    , 24'd4325    , 24'd4336    , 
//     24'd4346    , 24'd4357    , 24'd4367    , 24'd4378    , 24'd4388    , 24'd4398    , 24'd4409    , 24'd4419    , 
//     24'd4429    , 24'd4440    , 24'd4450    , 24'd4460    , 24'd4471    , 24'd4481    , 24'd4491    , 24'd4502    , 
//     24'd4512    , 24'd4522    , 24'd4533    , 24'd4543    , 24'd4553    , 24'd4564    , 24'd4574    , 24'd4584    , 
//     24'd4594    , 24'd4605    , 24'd4615    , 24'd4625    , 24'd4635    , 24'd4645    , 24'd4656    , 24'd4666    , 
//     24'd4676    , 24'd4686    , 24'd4696    , 24'd4707    , 24'd4717    , 24'd4727    , 24'd4737    , 24'd4747    , 
//     24'd4757    , 24'd4767    , 24'd4778    , 24'd4788    , 24'd4798    , 24'd4808    , 24'd4818    , 24'd4828    , 
//     24'd4838    , 24'd4848    , 24'd4858    , 24'd4868    , 24'd4878    , 24'd4888    , 24'd4898    , 24'd4909    , 
//     24'd4919    , 24'd4929    , 24'd4939    , 24'd4949    , 24'd4959    , 24'd4969    , 24'd4979    , 24'd4988    , 
//     24'd4998    , 24'd5008    , 24'd5018    , 24'd5028    , 24'd5038    , 24'd5048    , 24'd5058    , 24'd5068    , 
//     24'd5078    , 24'd5088    , 24'd5098    , 24'd5108    , 24'd5118    , 24'd5127    , 24'd5137    , 24'd5147    , 
//     24'd5157    , 24'd5167    , 24'd5177    , 24'd5187    , 24'd5196    , 24'd5206    , 24'd5216    , 24'd5226    , 
//     24'd5236    , 24'd5245    , 24'd5255    , 24'd5265    , 24'd5275    , 24'd5285    , 24'd5294    , 24'd5304    , 
//     24'd5314    , 24'd5324    , 24'd5333    , 24'd5343    , 24'd5353    , 24'd5362    , 24'd5372    , 24'd5382    , 
//     24'd5392    , 24'd5401    , 24'd5411    , 24'd5421    , 24'd5430    , 24'd5440    , 24'd5450    , 24'd5459    , 
//     24'd5469    , 24'd5479    , 24'd5488    , 24'd5498    , 24'd5507    , 24'd5517    , 24'd5527    , 24'd5536    , 
//     24'd5546    , 24'd5555    , 24'd5565    , 24'd5575    , 24'd5584    , 24'd5594    , 24'd5603    , 24'd5613    , 
//     24'd5622    , 24'd5632    , 24'd5641    , 24'd5651    , 24'd5661    , 24'd5670    , 24'd5680    , 24'd5689    , 
//     24'd5699    , 24'd5708    , 24'd5718    , 24'd5727    , 24'd5736    , 24'd5746    , 24'd5755    , 24'd5765    , 
//     24'd5774    , 24'd5784    , 24'd5793    , 24'd5803    , 24'd5812    , 24'd5821    , 24'd5831    , 24'd5840    , 
//     24'd5850    , 24'd5859    , 24'd5868    , 24'd5878    , 24'd5887    , 24'd5897    , 24'd5906    , 24'd5915    , 
//     24'd5925    , 24'd5934    , 24'd5943    , 24'd5953    , 24'd5962    , 24'd5971    , 24'd5981    , 24'd5990    , 
//     24'd5999    , 24'd6008    , 24'd6018    , 24'd6027    , 24'd6036    , 24'd6046    , 24'd6055    , 24'd6064    , 
//     24'd6073    , 24'd6083    , 24'd6092    , 24'd6101    , 24'd6110    , 24'd6119    , 24'd6129    , 24'd6138    , 
//     24'd6147    , 24'd6156    , 24'd6165    , 24'd6175    , 24'd6184    , 24'd6193    , 24'd6202    , 24'd6211    , 
//     24'd6221    , 24'd6230    , 24'd6239    , 24'd6248    , 24'd6257    , 24'd6266    , 24'd6275    , 24'd6284    , 
//     24'd6294    , 24'd6303    , 24'd6312    , 24'd6321    , 24'd6330    , 24'd6339    , 24'd6348    , 24'd6357    , 
//     24'd6366    , 24'd6375    , 24'd6384    , 24'd6393    , 24'd6402    , 24'd6411    , 24'd6421    , 24'd6430    , 
//     24'd6439    , 24'd6448    , 24'd6457    , 24'd6466    , 24'd6475    , 24'd6484    , 24'd6493    , 24'd6502    , 
//     24'd6511    , 24'd6519    , 24'd6528    , 24'd6537    , 24'd6546    , 24'd6555    , 24'd6564    , 24'd6573    , 
//     24'd6582    , 24'd6591    , 24'd6600    , 24'd6609    , 24'd6618    , 24'd6627    , 24'd6636    , 24'd6644    , 
//     24'd6653    , 24'd6662    , 24'd6671    , 24'd6680    , 24'd6689    , 24'd6698    , 24'd6707    , 24'd6715    , 
//     24'd6724    , 24'd6733    , 24'd6742    , 24'd6751    , 24'd6760    , 24'd6768    , 24'd6777    , 24'd6786    , 
//     24'd6795    , 24'd6804    , 24'd6812    , 24'd6821    , 24'd6830    , 24'd6839    , 24'd6847    , 24'd6856    , 
//     24'd6865    , 24'd6874    , 24'd6883    , 24'd6891    , 24'd6900    , 24'd6909    , 24'd6917    , 24'd6926    , 
//     24'd6935    , 24'd6944    , 24'd6952    , 24'd6961    , 24'd6970    , 24'd6978    , 24'd6987    , 24'd6996    , 
//     24'd7004    , 24'd7013    , 24'd7022    , 24'd7030    , 24'd7039    , 24'd7048    , 24'd7056    , 24'd7065    , 
//     24'd7074    , 24'd7082    , 24'd7091    , 24'd7099    , 24'd7108    , 24'd7117    , 24'd7125    , 24'd7134    , 
//     24'd7142    , 24'd7151    , 24'd7160    , 24'd7168    , 24'd7177    , 24'd7185    , 24'd7194    , 24'd7202    , 
//     24'd7211    , 24'd7220    , 24'd7228    , 24'd7237    , 24'd7245    , 24'd7254    , 24'd7262    , 24'd7271    , 
//     24'd7279    , 24'd7288    , 24'd7296    , 24'd7305    , 24'd7313    , 24'd7322    , 24'd7330    , 24'd7339    , 
//     24'd7347    , 24'd7356    , 24'd7364    , 24'd7372    , 24'd7381    , 24'd7389    , 24'd7398    , 24'd7406    , 
//     24'd7415    , 24'd7423    , 24'd7432    , 24'd7440    , 24'd7448    , 24'd7457    , 24'd7465    , 24'd7474    , 
//     24'd7482    , 24'd7490    , 24'd7499    , 24'd7507    , 24'd7515    , 24'd7524    , 24'd7532    , 24'd7541    , 
//     24'd7549    , 24'd7557    , 24'd7566    , 24'd7574    , 24'd7582    , 24'd7591    , 24'd7599    , 24'd7607    , 
//     24'd7616    , 24'd7624    , 24'd7632    , 24'd7640    , 24'd7649    , 24'd7657    , 24'd7665    , 24'd7674    , 
//     24'd7682    , 24'd7690    , 24'd7698    , 24'd7707    , 24'd7715    , 24'd7723    , 24'd7731    , 24'd7740    , 
//     24'd7748    , 24'd7756    , 24'd7764    , 24'd7773    , 24'd7781    , 24'd7789    , 24'd7797    , 24'd7805    , 
//     24'd7814    , 24'd7822    , 24'd7830    , 24'd7838    , 24'd7846    , 24'd7855    , 24'd7863    , 24'd7871    , 
//     24'd7879    , 24'd7887    , 24'd7895    , 24'd7903    , 24'd7912    , 24'd7920    , 24'd7928    , 24'd7936    , 
//     24'd7944    , 24'd7952    , 24'd7960    , 24'd7969    , 24'd7977    , 24'd7985    , 24'd7993    , 24'd8001    , 
//     24'd8009    , 24'd8017    , 24'd8025    , 24'd8033    , 24'd8041    , 24'd8049    , 24'd8057    , 24'd8065    , 
//     24'd8074    , 24'd8082    , 24'd8090    , 24'd8098    , 24'd8106    , 24'd8114    , 24'd8122    , 24'd8130    , 
//     24'd8138    , 24'd8146    , 24'd8154    , 24'd8162    , 24'd8170    , 24'd8178    , 24'd8186    , 24'd8194    , 
//     24'd8202    , 24'd8210    , 24'd8218    , 24'd8226    , 24'd8234    , 24'd8242    , 24'd8250    , 24'd8258    , 
//     24'd8265    , 24'd8273    , 24'd8281    , 24'd8289    , 24'd8297    , 24'd8305    , 24'd8313    , 24'd8321    , 
//     24'd8329    , 24'd8337    , 24'd8345    , 24'd8353    , 24'd8361    , 24'd8368    , 24'd8376    , 24'd8384    , 
//     24'd8392    , 24'd8400    , 24'd8408    , 24'd8416    , 24'd8424    , 24'd8431    , 24'd8439    , 24'd8447    , 
//     24'd8455    , 24'd8463    , 24'd8471    , 24'd8478    , 24'd8486    , 24'd8494    , 24'd8502    , 24'd8510    , 
//     24'd8517    , 24'd8525    , 24'd8533    , 24'd8541    , 24'd8549    , 24'd8556    , 24'd8564    , 24'd8572    , 
//     24'd8580    , 24'd8588    , 24'd8595    , 24'd8603    , 24'd8611    , 24'd8619    , 24'd8626    , 24'd8634    , 
//     24'd8642    , 24'd8650    , 24'd8657    , 24'd8665    , 24'd8673    , 24'd8681    , 24'd8688    , 24'd8696    , 
//     24'd8704    , 24'd8711    , 24'd8719    , 24'd8727    , 24'd8734    , 24'd8742    , 24'd8750    , 24'd8757    , 
//     24'd8765    , 24'd8773    , 24'd8781    , 24'd8788    , 24'd8796    , 24'd8803    , 24'd8811    , 24'd8819    , 
//     24'd8826    , 24'd8834    , 24'd8842    , 24'd8849    , 24'd8857    , 24'd8865    , 24'd8872    , 24'd8880    , 
//     24'd8887    , 24'd8895    , 24'd8903    , 24'd8910    , 24'd8918    , 24'd8925    , 24'd8933    , 24'd8941    , 
//     24'd8948    , 24'd8956    , 24'd8963    , 24'd8971    , 24'd8978    , 24'd8986    , 24'd8994    , 24'd9001    , 
//     24'd9009    , 24'd9016    , 24'd9024    , 24'd9031    , 24'd9039    , 24'd9046    , 24'd9054    , 24'd9061    , 
//     24'd9069    , 24'd9076    , 24'd9084    , 24'd9091    , 24'd9099    , 24'd9106    , 24'd9114    , 24'd9121    , 
//     24'd9129    , 24'd9136    , 24'd9144    , 24'd9151    , 24'd9159    , 24'd9166    , 24'd9174    , 24'd9181    , 
//     24'd9189    , 24'd9196    , 24'd9204    , 24'd9211    , 24'd9218    , 24'd9226    , 24'd9233    , 24'd9241    , 
//     24'd9248    , 24'd9256    , 24'd9263    , 24'd9270    , 24'd9278    , 24'd9285    , 24'd9293    , 24'd9300    , 
//     24'd9307    , 24'd9315    , 24'd9322    , 24'd9330    , 24'd9337    , 24'd9344    , 24'd9352    , 24'd9359    , 
//     24'd9366    , 24'd9374    , 24'd9381    , 24'd9388    , 24'd9396    , 24'd9403    , 24'd9410    , 24'd9418    , 
//     24'd9425    , 24'd9432    , 24'd9440    , 24'd9447    , 24'd9454    , 24'd9462    , 24'd9469    , 24'd9476    , 
//     24'd9484    , 24'd9491    , 24'd9498    , 24'd9506    , 24'd9513    , 24'd9520    , 24'd9527    , 24'd9535    , 
//     24'd9542    , 24'd9549    , 24'd9556    , 24'd9564    , 24'd9571    , 24'd9578    , 24'd9586    , 24'd9593    , 
//     24'd9600    , 24'd9607    , 24'd9614    , 24'd9622    , 24'd9629    , 24'd9636    , 24'd9643    , 24'd9651    , 
//     24'd9658    , 24'd9665    , 24'd9672    , 24'd9679    , 24'd9687    , 24'd9694    , 24'd9701    , 24'd9708    , 
//     24'd9715    , 24'd9723    , 24'd9730    , 24'd9737    , 24'd9744    , 24'd9751    , 24'd9758    , 24'd9766    , 
//     24'd9773    , 24'd9780    , 24'd9787    , 24'd9794    , 24'd9801    , 24'd9809    , 24'd9816    , 24'd9823    , 
//     24'd9830    , 24'd9837    , 24'd9844    , 24'd9851    , 24'd9858    , 24'd9866    , 24'd9873    , 24'd9880    , 
//     24'd9887    , 24'd9894    , 24'd9901    , 24'd9908    , 24'd9915    , 24'd9922    , 24'd9929    , 24'd9936    , 
//     24'd9944    , 24'd9951    , 24'd9958    , 24'd9965    , 24'd9972    , 24'd9979    , 24'd9986    , 24'd9993    
// };