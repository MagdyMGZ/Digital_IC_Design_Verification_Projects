package sa_pkg;
localparam TESTS = 1000;
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "sa_config.svh"
`include "sa_sequence_item.svh"
`include "sa_sequencer.svh"
`include "sa_sequence.svh"
`include "sa_driver.svh"
`include "sa_monitor.svh"
`include "sa_agent.svh"
`include "sa_scoreboard.svh"
`include "sa_collector.svh"
`include "sa_env.svh"
`include "sa_test.svh"
endpackage